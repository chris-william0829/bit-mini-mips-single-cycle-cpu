//`timescale 1ns / 1ps
`include "ControlSignalDefine.v"
//////////////////////////////////////////////////////////////////////////////////
// Company: BIT
// Engineer: Chris
// 
// Create Date: 2021/08/26 16:18:49
// Design Name: NextPC
// Module Name: NextPC
// Project Name: single cycle mips cpu
// Target Devices: 
// Tool Versions: vivado 2019.2
// Description: select the next pc by the signal generated by instruction
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module NextPC(
    input [31:0] PC,
    input [2:0] NextPCSignal,
    input [25:0] JumpAddr,
    input [31:0] JumpReg,
    output reg[31:0] NextPC
    );
    wire [31:0] PC4;
    assign PC4 = PC + 4;
    always @ (*) begin
        case (NextPCSignal)
            `PC_PLUS4: NextPC <= PC4;
            `PC_BRANCH: NextPC <= PC4 + { {14{JumpAddr[15]}}, JumpAddr[15:0], 2'b00};   //Branch
            `PC_IMM: NextPC <= {PC4[31:28],JumpAddr[25:0],2'b00};       //j,jal
            `PC_REG: NextPC <= JumpReg;                                 //jr,jalr
            `PC_HALT: NextPC <= PC;                                     //halt
            default: NextPC <= `ZeroWord;
        endcase
    end
    
endmodule
